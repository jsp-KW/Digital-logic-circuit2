module cla4_ov(a,b,ci,s,c3,co);
	input [3:0] a,b; //4bit input signal a,b
	input ci;// 1bit input signal ci
	output[3:0] s;// 4bit output signal s
	output c3,co;// 1bit output signal c3,co
	
	wire c1, c2; //1bit wire c1,c2
	
	fa_v2 U0_fa (.a(a[0]),.b(b[0]),.ci(ci),.s(s[0])); //instance name U0_fa, use fa_v2 module
	fa_v2 U1_fa (.a(a[1]),.b(b[1]),.ci(c1),.s(s[1])); //instance name U1_fa, use fa_v2 module
	fa_v2 U2_fa (.a(a[2]),.b(b[2]),.ci(c2),.s(s[2])); //instance name U2_fa, use fa_v2 module
	fa_v2 U3_fa (.a(a[3]),.b(b[3]),.ci(c3),.s(s[3])); //instance name U3_fa, use fa_v2 module
	clb  U4_clb4(.a(a), .b(b), .ci(ci), .c1(c1), .c2(c2), .c3(c3), .co(co));  //instance name U4_clb4, use clb module

endmodule
