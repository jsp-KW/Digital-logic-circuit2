module mx2_4bits(d0,d1,s,y);
	
	input [3:0]d0, d1; // 4bit input signal d0, d1
	input s; // 1bit input signal s
	output [3:0]y; // 1bit output signal y
	
	//module instance, use mx2 module//
	mx2 mx2_U0(.d0(d0[0]), .d1(d1[0]), .s(s), .y(y[0])); 
	mx2 mx2_U1(.d0(d0[1]), .d1(d1[1]), .s(s), .y(y[1]));
	mx2 mx2_U2(.d0(d0[2]), .d1(d1[2]), .s(s), .y(y[2]));
	mx2 mx2_U3(.d0(d0[3]), .d1(d1[3]), .s(s), .y(y[3]));
	
endmodule
